//module load(input clk, data,
//	input [15:0] C,
//	output readEnable
//	);