module array_divider (
	input wire [6:0] a,
	input wire [3:0] b,
	input wire mode,
	output wire [3:0] q,
	output wire [3:0] r
);

	wire mode1, mode2, mode3, mode4;
	wire mode5, mode6, mode7, mode8;
	wire mode9, mode10, mode11, mode12;
	wire mode13, mode14, mode15, mode16;
	
endmodule